interface intf;
  
  logic d;
  logic q;
  logic reset;
  
endinterface
