interface intf#(parameter WIDTH = 4,ADDRESS = 4 );
  
  logic clk;
  logic reset;
  logic up;
  logic down;
  logic reset;
  logic [3:0]count;
  
  
endinterface
