interface intf();
  
  logic a;
  logic b;
  logic c;
  logic sum;
  logic carry;
  
  modport dut( input a,b,c , output sum,carry );
  
endinterface
